ENTITY Calculadora IS



END Calculadora;

architecture  of Calculadora is



begin





   
